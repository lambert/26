.TITLE OCTAVE FILTER - MAIN BOARD - INPUT STAGE - FREQUENCY RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 pulse(iv=0 pv=15 rise=.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=.01)

VS 1 0 AC 1 SIN(0 1 16k)
C1 1 2 680n
R1 0 2 100k
R2 2 6 10K
R3 3 7 47k
R4 7 0 4700
XOP1 6 7 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT TRAN V(1) V(3)

*     FROM  TO    STEP
.TRAN 0     0.01  0.000001 TRACE ALL

.END
