.TITLE OCTAVE FILTER - FUNCTION 018: 8 KHZ BAND-PASS FILTER - TRANSIENT RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 pulse(iv=0 pv=15 rise=0.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=0.01)

VS 1 0 AC 1 SIN(0 1.41 31.5)
R1 1 2 26.7k
R2 3 6 267K
R3 0 2 14700
C1 2 6 470pF
C2 3 2 470pF
XOP1 0 6 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT TRAN V(1) V(3) V(4) V(5)

*     FROM  TO   STEP
.TRAN 0     0.1  0.00001 TRACE ALL

.END
