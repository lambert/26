.TITLE OCTAVE FILTER - FUNCTION 012: 1 kHZ BAND-PASS FILTER - FREQUENCY RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 15
VEE 5 0 -15

VS 1 0 AC 1 SIN(0 1.41 1k)
R1 1 2 21.3k
R2 3 6 213K
R3 0 2 8300
C1 2 6 4.7nF
C2 3 2 4.7nF
XOP1 0 6 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT AC VDB(3)

*     FROM      TO   STEP
.TRAN 0.00001   0.2  0.0001

*       #STEPS/DECADE FROM   TO 
.AC DEC 20            0.1    100k

.END
