.TITLE OCTAVE FILTER - MAIN BOARD - INPUT STAGE - FREQUENCY RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 15
VEE 5 0 -15

VS 1 0 AC 1 SIN(0 0.1 100)
C1 1 2 680n
R1 0 2 100k
R2 2 6 10K
R3 3 7 47k
R4 7 0 4700
XOP1 6 7 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT AC VDB(3)

*     FROM      TO   STEP
.TRAN 0.00001   0.2  0.0001

*       #STEPS/DECADE FROM   TO 
.AC DEC 20            0.01   10Meg

.END
