.TITLE OCTAVE FILTER - FUNCTION 007: 125 HZ DETECTOR - TRANSIENT RESPONSE

.INCLUDE UA741.subckt

.MODEL 1N4148 D IS=2e-14


VCC 4 0 pulse(iv=0 pv=15 rise=0.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=0.01)

VS 1 0 AC 1 SIN(0 1.41 125)
C1 0 7 1uF
D1 2 3 1N4148
D2 3 6 1N4148
R1 1 2 10000
R2 6 7 1000
R3 8 2 15000
R4 0 9 10000
R5 8 9 .001
XOP1 0 2 0 4 5 3 UA741
XOP2 7 8 0 4 5 9 UA741


.PRINT OP Iter(0) V(3)

.PRINT TRAN I(R1) I(R2) I(R3) I(R4) I(R5) I(D1) I(D2)

*     FROM  TO   STEP
.TRAN 0     0.1  0.00001

.END
