.TITLE OCTAVE FILTER - FUNCTION 018: 8 kHZ BAND-PASS FILTER - FREQUENCY RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 15
VEE 5 0 -15

VS 1 0 AC 1 SIN(0 1.41 8k)
R1 1 2 26.7k
R2 3 6 267K
R3 0 2 14700
C1 2 6 470pF
C2 3 2 470pF
XOP1 0 6 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT AC VDB(3)

*     FROM      TO   STEP
.TRAN 0.00001   0.2  0.0001

*       #STEPS/DECADE FROM   TO 
.AC DEC 20            0.1    100k

.END
