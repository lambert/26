.TITLE OCTAVE FILTER - 31.5 HZ MODULE - SECOND STAGE - TRANSIENT RESPONSE

VCC 4 0 pulse(iv=0 pv=15 rise=.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=.01)

.MODEL 1N4148 D IS=2e-14

VS 1 0 AC 1 SIN(0 4.138 31.5)
C1 0 7 1uF
D1 2 3 1N4148
D2 3 6 1N4148
R1 1 2 10000
R2 6 7 1000
R3 8 2 15000
R4 0 9 10000
R5 8 9 .001
XOP1 0 2 0 4 5 3 UA741
XOP2 7 8 0 4 5 9 UA741

.SUBCKT UA741    1   2   3   4    5    6
*               Vi+ Vi- GND PWR+ PWR- Vout
Q1 11 1 13 OPNPN1
Q2 12 2 14 OPNPN2
RC1 4 11 5.305165E+03
RC2 4 12 5.305165E+03
C1 11 12 5.459553E-12
RE1 13 10 2.151297E+03
RE2 14 10 2.151297E+03
IEE 10 5 1.666000E-05
CE  10 3 3.000000E-12
RE  10 3 1.200480E+07
GCM 3 21 10 3 5.960753E-09
GA 21 3 12 11 1.884955E-04
R2 21 3 1.000000E+05
C2 21 22 3.000000E-11
GB 22 3 21 3 2.357851E+02
RO2 22 3 4.500000E+01
D1 22 31 OPD12
D2 31 22 OPD12
EC 31 3 6 3 1.0
RO1 22 6 3.000000E+01
D3 6 24 OPD34
VC 4 24 2.803238E+00
D4 25 6 OPD34
VE 25 5 2.803238E+00
.MODEL OPD12 D (IS=9.762287E-11)
.MODEL OPD34 D (IS=8.000000E-16)
.MODEL OPNPN1 NPN (IS=8.000000E-16 BF=9.166667E+01)
.MODEL OPNPN2 NPN (IS=8.309478E-16 BF=1.178571E+02)
.ENDS


.PRINT OP Iter(0) V(3)

.PRINT TRAN V(1) V(3) V(9)

*     FROM  TO   STEP
.TRAN 0.2   0.3  0.00001

.END
