.TITLE OCTAVE FILTER - FUNCTION 004: 63 HZ BAND-PASS FILTER - TRANSIENT RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 pulse(iv=0 pv=15 rise=0.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=0.01)

VS 1 0 AC 1 SIN(0 1.41 16k)
R1 1 2 15900
R2 3 6 159K
R3 0 2 7200
C1 2 6 100nF
C2 3 2 100nF
XOP1 0 6 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT TRAN V(1) V(3) V(4) V(5)

*     FROM  TO   STEP
.TRAN 0     0.1  0.00001 TRACE ALL

.END
