.TITLE OCTAVE FILTER - FUNCTION 020: 16 KHZ BAND-PASS FILTER - TRANSIENT RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 pulse(iv=0 pv=15 rise=0.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=0.01)

VS 1 0 AC 1 SIN(0 1.41 16k)
R1 1 2 28k
R2 3 6 280K
R3 0 2 14700
C1 2 6 220pF
C2 3 2 220pF
XOP1 0 6 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT TRAN P(R1) P(R2) P(R3)

*     FROM  TO   STEP
.TRAN 0     0.02  0.00001 TRACE ALL

.END
