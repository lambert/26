.TITLE OCTAVE FILTER - FUNCTION 004: 63 HZ BAND-PASS FILTER - TRANSIENT RESPONSE

.INCLUDE UA741.subckt


VCC 4 0 pulse(iv=0 pv=15 rise=0.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=0.01)

VS 1 0 AC 1 SIN(0 1.41 63)
R1 1 2 15900
R2 3 6 159K
R3 0 2 7200
C1 2 6 100nF
C2 3 2 100nF
XOP1 0 6 0 4 5 3 UA741


.PRINT OP Iter(0) V(3)

.PRINT TRAN I(R1) I(R2) I(R3)

*     FROM  TO   STEP
.TRAN 0     0.2  0.0001 TRACE ALL

.END
