.TITLE OCTAVE FILTER - FIRST STAGE - TRANSIENT RESPONSE

VCC 4 0 pulse(iv=0 pv=15 rise=.01)
VEE 5 0 pulse(iv=0 pv=-15 rise=.01)

VS 1 0 AC 1 SIN(0 1 31.5)
R1 1 2 14200
R2 3 6 142K
R3 0 2 7200
C1 2 6 220nF
C2 3 2 220nF
XOP1 0 6 4 5 3 CA3140


*$ model description: "awbca3140"
*a Device model created by analog_uprev for ca3140 on Thu Mar 1 18:48:14 IST 2001
* CONNECTIONS:   NON-INVERTING INPUT
*                |  INVERTING INPUT
*                |  |  POSITIVE POWER SUPPLY
*                |  |  |  NEGATIVE POWER SUPPLY
*                |  |  |  |  OUTPUT
*                |  |  |  |  |
.subckt CA3140   1  36 15 20 12
*START OF DECK
* +IN -IN OUT +VSS -VSS
*NODE: 1 36 15 20 12
*------INPUT STAGE-------
VOSBAL 7 29 3.00000000E-03
EU1 8 1 20 12 0.0001
EU2 8 7 5 12 -1
*RB1 12 10 1 TC= 1.991040E-03 (-1.244400E-04)
IB4 10 12 1.000000E-06
*RB3 12 5 8743.17 TC= 1.60000000E-03 (0.00000000E+00)
IB3 12 5 5.718750E-07
G1 12 1 10 12 1.025000E-05
G2 12 36 10 12 9.750000E-06
RDM 36 29 1.500000E+12
RCM 31 13 1.500000E+12
CDM 36 29 4.000000E-12
G5 31 13 36 31 6.66667E-13
G6 31 13 1 31 6.66667E-13
*------INTERMEDIATE STAGE-------
GDM 31 16 29 36 1
GCM 31 16 13 31 -1.58113883E-05
R1 31 16 3.16358380E+02
C1 31 16 6.45457E-11
VCP 23 31 100
VCM 24 31 -100
DD1 16 23 MD2
.MODEL MD2 D XTI=1.000000P
* SPECTRE: + IMAX=1000
DD2 24 16 MD2
G3 31 6 16 31 -1.07249255E-06
R2 31 6 100000
C2 11 6 1.2E-11
RP1 31 20 3750
RP2 31 12 3750
*------OUTPUT STAGE-------
G4 31 11 6 31 -5.10867719E+01
ROUT 31 11 60
DD3 11 9 MD3
.MODEL MD3 D IS=10.0F XTI=1.0P N= 3.612647E-01
* SPECTRE: + IMAX=1000
DD4 9 11 MD4
.MODEL MD4 D IS=10.0F XTI=1.0P N= 8.028126E-01
* SPECTRE: + IMAX=1000
EU6 9 31 2 31 1
RO1 11 26 20
FF1 31 28 VFF1 1
VFF1 26 2 0.0
FF2 31 20 VFF2 -1
VFF2 33 31 0.0
FF3 12 31 VFF3 -1
VFF3 31 27 0.0
DD8 27 28 MID
DD7 28 33 MID
.MODEL MID D XTI=1.000000F N=1 IS=10.000000F
* SPECTRE: + IMAX=1000
VP 20 22 -29.2613
VM 21 12 -29.3113
DD5 25 22 MID
DD6 21 17 MID
VP1 20 30 2.7501
VM1 32 12 .859456
DD9 2 30 MD9
DD10 32 15 MD9
.MODEL MD9 D XTI=1.000000F N=1 IS=10.000000F
* SPECTRE: + IMAX=1000
*HH1 25 2 POLY(2) VIC2 VIC1 0 1960 0 1540 0 0 0 0 0 0
*HH2 2 17 POLY(2) VIC3 VIC1 0 -1960 0 -1540 0 0 0 0 0 0
VIC1 37 3 0.0
VIC2 2 14 0.0
VIC3 14 15 0.0
VPP 37 0 1
RPP 3 0 100.0K
RO3 15 20 200.0MEG
RO2 15 12 200.0MEG
.ENDS
*$ end model description: "awbca3140"


.PRINT OP Iter(0) V(3)

.PRINT TRAN V(1) V(3)

*     FROM      TO   STEP
.TRAN 0.00001S  0.2S 0.0001S

.END
